module uart ();
input wire xmit_dataH_0, xmit_dataH_1, xmit_dataH_2, xmit_dataH_3, xmit_dataH_4, xmit_dataH_5, xmit_dataH_6, xmit_dataH_7, sys_clk, sys_rst_l, xmitH, uart_REC_dataH, test_mode, test_se, test_si;
output wire rec_dataH_0, rec_dataH_1, rec_dataH_2, rec_dataH_3, rec_dataH_4, rec_dataH_5, rec_dataH_6, rec_dataH_7, uart_XMIT_dataH, xmit_doneH, rec_readyH, test_so;
  assign test_pointTM  = test_mode;
  assign test_so = rec_dataH_temp[7];
  AND2X4 U305 (iCTRL, iXMIT_state_1_temp, iXMIT_state_1_);
  AND2X4 U303 (iCTRL, xmit_doneH_temp, xmit_doneH);
  ISOLORX8 U302 (iXMIT_CRTL, iRECEIVER_CTRL, iCTRL);
  OR4X4 U301 (iRECEIVER_state_CTRL, iRECEIVER_N_CTRL_1_, iRECEIVER_N_CTRL_2_, iRECEIVER_bitCell_CTRL, iRECEIVER_CTRL);
  NAND4X1 U300 (iRECEIVER_N18, iRECEIVER_N17, iRECEIVER_bitCell_cntrH_0_, iRECEIVER_bitCell_cntrH_1_, iRECEIVER_bitCell_CTRL);
  NAND4X1 U299 (iRECEIVER_N22, iRECEIVER_N21, iRECEIVER_N20, iRECEIVER_N19, iRECEIVER_N_CTRL_2_);
  NAND4X1 U298 (iRECEIVER_N28, iRECEIVER_N27, iRECEIVER_N26, iRECEIVER_N23, iRECEIVER_N_CTRL_1_);
  NAND4X1 U297 (iRECEIVER_next_state_2_, iRECEIVER_state_0_, iRECEIVER_state_1_, iRECEIVER_state_2_, iRECEIVER_state_CTRL);
  OR4X4 U296 (1'b0, iXMIT_N_CTRL_1_, iXMIT_N_CTRL_2_, iXMIT_xmit_CTRL, iXMIT_CRTL);
  NAND4X1 U295 (iXMIT_N24, iXMIT_xmit_ShiftRegH_7_, iXMIT_xmit_ShiftRegH_6_, iXMIT_xmit_ShiftRegH_5_, iXMIT_xmit_CTRL);
  NAND4X1 U294 (iXMIT_N28, iXMIT_N27, iXMIT_N26, iXMIT_N25, iXMIT_N_CTRL_2_);
  NAND4X1 U293 (n251, n239, n242, n246, iXMIT_N_CTRL_1_);
  XOR2X2 U230 (iRECEIVER_recd_bitCntrH_3_, n275, iRECEIVER_N28);
  NOR2X4 U229 (n274, n250, n275);
  XOR2X2 U228 (n250, n274, iRECEIVER_N27);
  XOR2X2 U227 (iRECEIVER_recd_bitCntrH_1_, iRECEIVER_recd_bitCntrH_0_, iRECEIVER_N26);
  XOR2X2 U226 (iRECEIVER_bitCell_cntrH_3_, n273, iRECEIVER_N19);
  NOR2X4 U225 (n272, n249, n273);
  XOR2X2 U224 (n249, n272, iRECEIVER_N18);
  XOR2X2 U223 (iRECEIVER_bitCell_cntrH_1_, iRECEIVER_bitCell_cntrH_0_, iRECEIVER_N17);
  XOR2X2 U222 (iXMIT_bitCountH_3_, n271, iXMIT_N46);
  NOR2X4 U221 (n270, n247, n271);
  XOR2X2 U220 (n247, n270, iXMIT_N45);
  XOR2X2 U219 (iXMIT_bitCountH_1_, iXMIT_bitCountH_0_, iXMIT_N44);
  XOR2X2 U218 (iXMIT_bitCell_cntrH_3_, n269, iXMIT_N25);
  NOR2X4 U217 (n268, n251, n269);
  XOR2X2 U216 (n251, n268, iXMIT_N24);
  XOR2X2 U215 (iXMIT_bitCell_cntrH_1_, iXMIT_bitCell_cntrH_0_, iXMIT_N23);
  INVX32 U214 (n64, n28);
  NAND2X4 U213 (n55, n56, iXMIT_xmit_doneInH);
  NAND2X4 U212 (iRECEIVER_bitCell_cntrH_1_, iRECEIVER_bitCell_cntrH_0_, n272);
  NAND2X4 U211 (iXMIT_bitCell_cntrH_1_, iXMIT_bitCell_cntrH_0_, n268);
  NAND2X4 U210 (iRECEIVER_recd_bitCntrH_1_, iRECEIVER_recd_bitCntrH_0_, n274);
  NAND2X4 U209 (n61, n69, n53);
  NAND2X4 U208 (iXMIT_bitCountH_1_, iXMIT_bitCountH_0_, n270);
  NAND2X4 U207 (n63, n44, iXMIT_next_state_1_);
  NAND2X4 U206 (xmit_dataH[7], n26, n43);
  NAND2X4 U205 (n42, n43, n211);
  NAND2X4 U204 (n67, n68, iXMIT_next_state_0_);
  INVX32 U202 (n8, n18);
  NAND2X4 U201 (n80, n91, n83);
  NAND4X1 U138 (iRECEIVER_bitCell_cntrH_3_, iRECEIVER_bitCell_cntrH_2_, iRECEIVER_bitCell_cntrH_1_, n255, n91);
  INVX32 U137 (n91, n79);
  AOI21X2 U135 (n79, iRECEIVER_state_0_, n241, n93);
  NAND4X1 U132 (iRECEIVER_bitCell_cntrH_2_, n255, n244, n256, n85);
  INVX32 U131 (n85, n88);
  AOI21X2 U129 (n88, n245, iRECEIVER_state_2_, n94);
  AND2X4 U128 (n93, n94, n92);
  AND2X4 U127 (n255, n92, iRECEIVER_N20);
  AND2X4 U126 (iRECEIVER_N17, n92, iRECEIVER_N21);
  AND2X4 U125 (iRECEIVER_N18, n92, iRECEIVER_N22);
  AND2X4 U124 (iRECEIVER_N19, n92, iRECEIVER_N23);
  NOR2X4 U123 (n241, n245, n80);
  NOR2X4 U120 (iRECEIVER_recd_bitCntrH_2_, iRECEIVER_recd_bitCntrH_1_, n89);
  NAND4X1 U118 (n80, iRECEIVER_recd_bitCntrH_3_, n89, n243, n86);
  AOI22X2 U117 (n88, iRECEIVER_state_1_, iRECEIVER_rec_datH, n241, n87);
  NAND4X1 U116 (n83, n238, n86, n87, iRECEIVER_next_state_0_);
  AOI21X2 U114 (iRECEIVER_state_1_, n85, n248, n84);
  ISOLORX8 U113 (iRECEIVER_state_0_, n84, n81);
  NAND3X4 U112 (n241, n238, n248, n82);
  NOR2X4 U111 (n238, iRECEIVER_state_0_, n8);
  NAND4X1 U109 (n81, n82, n18, n83, iRECEIVER_next_state_1_);
  AND2X4 U108 (n79, n80, iRECEIVER_next_state_2_);
  NAND3X4 U107 (n241, n238, iRECEIVER_rec_datH, n77);
  OAI21X2 U106 (n238, n245, n77, iRECEIVER_rec_readyInH);
  NAND3X4 U102 (iXMIT_bitCell_cntrH_2_, iXMIT_bitCell_cntrH_1_, iXMIT_bitCell_cntrH_3_, n75);
  NOR2X4 U101 (n254, n75, n57);
  NOR2X4 U100 (n242, n57, n62);
  INVX32 U99 (n62, n72);
  NOR2X4 U97 (n246, iXMIT_state_0_, n66);
  INVX32 U96 (n57, n74);
  NOR2X4 U95 (n246, n239, n54);
  NOR2X4 U94 (n75, iXMIT_bitCell_cntrH_0_, n61);
  INVX32 U93 (n61, n65);
  AOI22X2 U92 (n66, n74, n54, n65, n73);
  OAI21X2 U91 (n239, n72, n73, n71);
  AND2X4 U90 (n254, n71, iXMIT_N26);
  AND2X4 U89 (iXMIT_N23, n71, iXMIT_N27);
  AND2X4 U88 (iXMIT_N24, n71, iXMIT_N28);
  AND2X4 U87 (iXMIT_N25, n71, iXMIT_N29);
  OR4X4 U85 (n253, iXMIT_bitCountH_0_, iXMIT_bitCountH_1_, iXMIT_bitCountH_2_, n69);
  AOI22X2 U83 (n54, n53, iXMIT_state_2_, n239, n67);
  AOI21X2 U82 (n66, n57, n62, n68);
  AOI21X2 U80 (iXMIT_state_1_temp, n65, n66, n63);
  NAND3X4 U79 (n246, n242, xmitH, n64);
  AOI21X2 U77 (n239, iXMIT_state_2_, n28, n44);
  AOI22X2 U75 (n54, n61, n62, iXMIT_state_0_, n60);
  INVX32 U74 (n60, iXMIT_next_state_2_);
  INVX32 U73 (xmitH, n58);
  NAND3X4 U72 (n242, n58, n246, n55);
  NAND3X4 U71 (iXMIT_state_2_, iXMIT_state_0_, n57, n56);
  INVX32 U69 (n55, n51);
  INVX32 U68 (n54, n52);
  NOR2X4 U67 (n52, n53, n47);
  NOR2X4 U66 (n51, n47, n46);
  AOI22X2 U65 (iXMIT_bitCountH_0_, n46, n252, n47, n50);
  INVX32 U64 (n50, n223);
  AOI22X2 U63 (iXMIT_bitCountH_1_, n46, iXMIT_N44, n47, n49);
  INVX32 U62 (n49, n220);
  AOI22X2 U61 (iXMIT_bitCountH_2_, n46, iXMIT_N45, n47, n48);
  INVX32 U60 (n48, n217);
  AOI22X2 U59 (n46, iXMIT_bitCountH_3_, iXMIT_N46, n47, n45);
  INVX32 U58 (n45, n214);
  NOR2X4 U57 (n44, n28, n29);
  AOI21X2 U56 (iXMIT_xmit_ShiftRegH_7_, n44, n29, n42);
  INVX32 U55 (n44, n26);
  AOI22X2 U51 (xmit_dataH[6], n28, iXMIT_xmit_ShiftRegH_7_, n29, n41);
  OAI21X2 U50 (n26, n258, n41, n208);
  AOI22X2 U48 (xmit_dataH[5], n28, iXMIT_xmit_ShiftRegH_6_, n29, n39);
  OAI21X2 U47 (n26, n259, n39, n205);
  AOI22X2 U45 (xmit_dataH[4], n28, iXMIT_xmit_ShiftRegH_5_, n29, n37);
  OAI21X2 U44 (n26, n260, n37, n202);
  AOI22X2 U42 (xmit_dataH[3], n28, iXMIT_xmit_ShiftRegH_4_, n29, n35);
  OAI21X2 U41 (n26, n261, n35, n199);
  AOI22X2 U39 (xmit_dataH[2], n28, iXMIT_xmit_ShiftRegH_3_, n29, n33);
  OAI21X2 U38 (n26, n262, n33, n196);
  AOI22X2 U36 (xmit_dataH[1], n28, iXMIT_xmit_ShiftRegH_2_, n29, n31);
  OAI21X2 U35 (n263, n26, n31, n193);
  AOI22X2 U33 (xmit_dataH[0], n28, iXMIT_xmit_ShiftRegH_1_, n29, n27);
  OAI21X2 U32 (n257, n26, n27, n190);
  AOI22X2 U31 (iRECEIVER_rec_datH, n8, rec_dataH_rec[7], n18, n25);
  INVX32 U30 (n25, n165);
  AOI22X2 U29 (rec_dataH_rec[7], n8, rec_dataH_rec[6], n18, n24);
  INVX32 U28 (n24, n158);
  AOI22X2 U27 (rec_dataH_rec[6], n8, rec_dataH_rec[5], n18, n23);
  INVX32 U26 (n23, n151);
  AOI22X2 U25 (rec_dataH_rec[5], n8, rec_dataH_rec[4], n18, n22);
  INVX32 U24 (n22, n144);
  AOI22X2 U23 (rec_dataH_rec[4], n8, rec_dataH_rec[3], n18, n21);
  INVX32 U22 (n21, n137);
  AOI22X2 U21 (rec_dataH_rec[3], n8, rec_dataH_rec[2], n18, n20);
  INVX32 U20 (n20, n130);
  AOI22X2 U19 (rec_dataH_rec[2], n8, rec_dataH_rec[1], n18, n19);
  INVX32 U18 (n19, n123);
  AOI22X2 U17 (rec_dataH_rec[1], n8, rec_dataH_rec_0_temp, n18, n17);
  INVX32 U16 (n17, n116);
  OAI21X2 U15 (iRECEIVER_state_1_, n248, n238, n15);
  OAI21X2 U14 (n238, n245, n15, n9);
  AOI22X2 U13 (iRECEIVER_N28, n8, iRECEIVER_recd_bitCntrH_3_, n9, n12);
  INVX32 U12 (n12, n109);
  AOI22X2 U11 (n243, n8, iRECEIVER_recd_bitCntrH_0_, n9, n11);
  INVX32 U10 (n11, n106);
  AOI22X2 U9 (iRECEIVER_N26, n8, iRECEIVER_recd_bitCntrH_1_, n9, n10);
  INVX32 U8 (n10, n103);
  AOI22X2 U7 (iRECEIVER_N27, n8, iRECEIVER_recd_bitCntrH_2_, n9, n7);
  INVX32 U6 (n7, n100);
  AOI21X2 U5 (n242, n239, n257, n3);
  AOI21X2 U4 (iXMIT_state_2_, iXMIT_state_0_, n3, n2);
  OAI21X2 U3 (iXMIT_state_2_, iXMIT_state_1_, n2, uart_XMIT_dataH);
  INVX32 U290 (n370, n371);
  NAND2X4 U289 (1'b1, test_pointTM, n370);
  DFFARX1 iXMIT_bitCell_cntrH_reg_2_ (n180, sys_clk, sys_rst_l, iXMIT_bitCell_cntrH_2_, n251);
  DFFARX1 iXMIT_state_reg_0_ (n179, sys_clk, sys_rst_l, iXMIT_state_0_, n239);
  DFFARX1 iXMIT_state_reg_2_ (n178, sys_clk, sys_rst_l, iXMIT_state_2_, n242);
  DFFARX1 iXMIT_state_reg_1_ (n177, sys_clk, sys_rst_l, iXMIT_state_1_temp, n246);
  DFFARX1 iXMIT_bitCountH_reg_0_ (n176, sys_clk, sys_rst_l, iXMIT_bitCountH_0_, n252);
  DFFARX1 iXMIT_bitCountH_reg_1_ (n175, sys_clk, sys_rst_l, iXMIT_bitCountH_1_);
  DFFARX1 iXMIT_bitCountH_reg_2_ (n174, sys_clk, sys_rst_l, iXMIT_bitCountH_2_, n247);
  DFFARX1 iXMIT_bitCountH_reg_3_ (n173, sys_clk, sys_rst_l, iXMIT_bitCountH_3_, n253);
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_7_ (n172, sys_clk, sys_rst_l, iXMIT_xmit_ShiftRegH_7_);
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_6_ (n171, sys_clk, sys_rst_l, iXMIT_xmit_ShiftRegH_6_, n258);
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_5_ (n170, sys_clk, sys_rst_l, iXMIT_xmit_ShiftRegH_5_, n259);
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_4_ (n169, sys_clk, sys_rst_l, iXMIT_xmit_ShiftRegH_4_, n260);
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_3_ (n168, sys_clk, sys_rst_l, iXMIT_xmit_ShiftRegH_3_, n261);
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_2_ (n167, sys_clk, sys_rst_l, iXMIT_xmit_ShiftRegH_2_, n262);
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_1_ (n166, sys_clk, sys_rst_l, iXMIT_xmit_ShiftRegH_1_, n263);
  DFFARX1 iXMIT_xmit_doneH_reg (n164, sys_clk, sys_rst_l, xmit_doneH_temp);
  DFFARX1 iRECEIVER_state_reg_1_ (n163, sys_clk, sys_rst_l, iRECEIVER_state_1_, n241);
  DFFASX1 iRECEIVER_state_reg_0_ (n162, sys_clk, sys_rst_l, iRECEIVER_state_0_, n245);
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_0_ (n161, sys_clk, sys_rst_l, iRECEIVER_bitCell_cntrH_0_, n255);
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_1_ (n160, sys_clk, sys_rst_l, iRECEIVER_bitCell_cntrH_1_, n244);
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_2_ (n159, sys_clk, sys_rst_l, iRECEIVER_bitCell_cntrH_2_, n249);
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_3_ (n157, sys_clk, sys_rst_l, iRECEIVER_bitCell_cntrH_3_, n256);
  DFFARX1 iRECEIVER_state_reg_2_ (n156, sys_clk, sys_rst_l, iRECEIVER_state_2_, n238);
  DFFARX1 iRECEIVER_rec_readyH_reg (n155, sys_clk, sys_rst_l, rec_readyH);
  DFFARX1 iRECEIVER_par_dataH_reg_7_ (n154, sys_clk, sys_rst_l, rec_dataH_rec[7]);
  DFFARX1 rec_dataH_temp_reg_7_ (n153, test_pointDOUT, sys_rst_l, rec_dataH_temp[7]);
  DFFARX1 rec_dataH_reg_7_ (n152, sys_clk, sys_rst_l, rec_dataH[7]);
  DFFARX1 iRECEIVER_par_dataH_reg_6_ (n150, sys_clk, sys_rst_l, rec_dataH_rec[6]);
  DFFARX1 rec_dataH_temp_reg_6_ (n149, test_pointDOUT, sys_rst_l, rec_dataH_temp[6]);
  DFFARX1 rec_dataH_reg_6_ (n148, sys_clk, sys_rst_l, rec_dataH[6]);
  DFFARX1 iRECEIVER_par_dataH_reg_5_ (n147, sys_clk, sys_rst_l, rec_dataH_rec[5]);
  DFFARX1 rec_dataH_temp_reg_5_ (n146, test_pointDOUT, sys_rst_l, rec_dataH_temp[5]);
  DFFARX1 rec_dataH_reg_5_ (n145, sys_clk, sys_rst_l, rec_dataH[5]);
  DFFARX1 iRECEIVER_par_dataH_reg_4_ (n143, sys_clk, sys_rst_l, rec_dataH_rec[4]);
  DFFARX1 rec_dataH_temp_reg_4_ (n142, test_pointDOUT, sys_rst_l, rec_dataH_temp[4]);
  DFFARX1 rec_dataH_reg_4_ (n141, sys_clk, sys_rst_l, rec_dataH[4]);
  DFFARX1 iRECEIVER_par_dataH_reg_3_ (n140, sys_clk, sys_rst_l, rec_dataH_rec[3]);
  DFFARX1 rec_dataH_temp_reg_3_ (n139, test_pointDOUT, sys_rst_l, rec_dataH_temp[3]);
  DFFARX1 rec_dataH_reg_3_ (n138, sys_clk, sys_rst_l, rec_dataH[3]);
  DFFARX1 iRECEIVER_par_dataH_reg_2_ (n136, sys_clk, sys_rst_l, rec_dataH_rec[2]);
  DFFARX1 rec_dataH_temp_reg_2_ (n135, test_pointDOUT, sys_rst_l, rec_dataH_temp[2]);
  DFFARX1 rec_dataH_reg_2_ (n134, sys_clk, sys_rst_l, rec_dataH[2]);
  DFFARX1 iRECEIVER_par_dataH_reg_1_ (n133, sys_clk, sys_rst_l, rec_dataH_rec[1]);
  DFFARX1 rec_dataH_temp_reg_1_ (n132, test_pointDOUT, sys_rst_l, rec_dataH_temp[1]);
  DFFARX1 rec_dataH_reg_1_ (n131, sys_clk, sys_rst_l, rec_dataH[1]);
  DFFARX1 iRECEIVER_par_dataH_reg_0_ (n129, sys_clk, sys_rst_l, rec_dataH_rec_0_temp);
  DFFARX1 rec_dataH_temp_reg_0_ (n128, test_pointDOUT, sys_rst_l, rec_dataH_temp[0]);
  DFFARX1 rec_dataH_reg_0_ (n127, sys_clk, sys_rst_l, rec_dataH[0]);
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_3_ (n126, sys_clk, sys_rst_l, iRECEIVER_recd_bitCntrH_3_);
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_0_ (n125, sys_clk, sys_rst_l, iRECEIVER_recd_bitCntrH_0_, n243);
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_1_ (n124, sys_clk, sys_rst_l, iRECEIVER_recd_bitCntrH_1_);
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_2_ (n122, sys_clk, sys_rst_l, iRECEIVER_recd_bitCntrH_2_, n250);
  DFFARX1 iXMIT_bitCell_cntrH_reg_3_ (n121, sys_clk, sys_rst_l, iXMIT_bitCell_cntrH_3_);
  DFFARX1 iXMIT_bitCell_cntrH_reg_0_ (n120, sys_clk, sys_rst_l, iXMIT_bitCell_cntrH_0_, n254);
  DFFARX1 iXMIT_bitCell_cntrH_reg_1_ (n119, sys_clk, sys_rst_l, iXMIT_bitCell_cntrH_1_);
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_0_ (n118, sys_clk, sys_rst_l, n281, n257);
  DFFASX1 iRECEIVER_rec_datSyncH_reg (n117, sys_clk, sys_rst_l, iRECEIVER_rec_datSyncH);
  DFFASX1 iRECEIVER_rec_datH_reg (n115, sys_clk, sys_rst_l, iRECEIVER_rec_datH, n248);
  MUX21X2 U291 (rec_readyH, sys_clk, n371, test_pointDOUT);
  MUX21X1 U1 (iRECEIVER_next_state_2_, iRECEIVER_state_1_, test_se, n156);
  MUX21X1 U2 (iRECEIVER_N23, iRECEIVER_bitCell_cntrH_2_, test_se, n157);
  MUX21X1 U34 (iRECEIVER_N22, iRECEIVER_bitCell_cntrH_1_, test_se, n159);
  MUX21X1 U37 (iRECEIVER_N21, iRECEIVER_bitCell_cntrH_0_, test_se, n160);
  MUX21X1 U40 (iRECEIVER_N20, test_si, test_se, n161);
  MUX21X1 U43 (iRECEIVER_next_state_0_, iRECEIVER_recd_bitCntrH_3_, test_se, n162);
  MUX21X1 U46 (iRECEIVER_next_state_1_, iRECEIVER_state_0_, test_se, n163);
  MUX21X1 U49 (iXMIT_xmit_doneInH, iXMIT_xmit_ShiftRegH_7_, test_se, n164);
  MUX21X1 U52 (n193, n281, test_se, n166);
  MUX21X1 U53 (n196, iXMIT_xmit_ShiftRegH_1_, test_se, n167);
  MUX21X1 U54 (n199, iXMIT_xmit_ShiftRegH_2_, test_se, n168);
  MUX21X1 U70 (n202, iXMIT_xmit_ShiftRegH_3_, test_se, n169);
  MUX21X1 U76 (n205, iXMIT_xmit_ShiftRegH_4_, test_se, n170);
  MUX21X1 U78 (n208, iXMIT_xmit_ShiftRegH_5_, test_se, n171);
  MUX21X1 U81 (n211, iXMIT_xmit_ShiftRegH_6_, test_se, n172);
  MUX21X1 U84 (n214, iXMIT_bitCountH_2_, test_se, n173);
  MUX21X1 U86 (n217, iXMIT_bitCountH_1_, test_se, n174);
  MUX21X1 U98 (n220, iXMIT_bitCountH_0_, test_se, n175);
  MUX21X1 U103 (n223, iXMIT_bitCell_cntrH_3_, test_se, n176);
  MUX21X1 U104 (iXMIT_next_state_1_, iXMIT_state_0_, test_se, n177);
  MUX21X1 U105 (iXMIT_next_state_2_, iXMIT_state_1_temp, test_se, n178);
  MUX21X1 U110 (iXMIT_next_state_0_, iXMIT_bitCountH_3_, test_se, n179);
  MUX21X1 U115 (iXMIT_N28, iXMIT_bitCell_cntrH_1_, test_se, n180);
  MUX21X1 U119 (iRECEIVER_rec_datSyncH, rec_dataH_rec[7], test_se, n115);
  MUX21X1 U121 (uart_REC_dataH, iRECEIVER_rec_datH, test_se, n117);
  MUX21X1 U122 (n190, iXMIT_state_2_, test_se, n118);
  MUX21X1 U130 (iXMIT_N27, iXMIT_bitCell_cntrH_0_, test_se, n119);
  MUX21X1 U133 (iXMIT_N26, iRECEIVER_state_2_, test_se, n120);
  MUX21X1 U134 (iXMIT_N29, iXMIT_bitCell_cntrH_2_, test_se, n121);
  MUX21X1 U136 (n100, iRECEIVER_recd_bitCntrH_1_, test_se, n122);
  MUX21X1 U139 (n103, iRECEIVER_recd_bitCntrH_0_, test_se, n124);
  MUX21X1 U140 (n106, rec_readyH, test_se, n125);
  MUX21X1 U141 (n109, iRECEIVER_recd_bitCntrH_2_, test_se, n126);
  MUX21X1 U142 (rec_dataH_temp[0], xmit_doneH_temp, test_se, n127);
  MUX21X1 U143 (rec_dataH_rec_0_temp, rec_dataH[7], test_se, n128);
  MUX21X1 U144 (n116, iRECEIVER_bitCell_cntrH_3_, test_se, n129);
  MUX21X1 U145 (rec_dataH_temp[1], rec_dataH[0], test_se, n131);
  MUX21X1 U146 (rec_dataH_rec[1], rec_dataH_temp[0], test_se, n132);
  MUX21X1 U147 (n123, rec_dataH_rec_0_temp, test_se, n133);
  MUX21X1 U148 (rec_dataH_temp[2], rec_dataH[1], test_se, n134);
  MUX21X1 U149 (rec_dataH_rec[2], rec_dataH_temp[1], test_se, n135);
  MUX21X1 U150 (n130, rec_dataH_rec[1], test_se, n136);
  MUX21X1 U151 (rec_dataH_temp[3], rec_dataH[2], test_se, n138);
  MUX21X1 U152 (rec_dataH_rec[3], rec_dataH_temp[2], test_se, n139);
  MUX21X1 U153 (n137, rec_dataH_rec[2], test_se, n140);
  MUX21X1 U154 (rec_dataH_temp[4], rec_dataH[3], test_se, n141);
  MUX21X1 U155 (rec_dataH_rec[4], rec_dataH_temp[3], test_se, n142);
  MUX21X1 U156 (n144, rec_dataH_rec[3], test_se, n143);
  MUX21X1 U157 (rec_dataH_temp[5], rec_dataH[4], test_se, n145);
  MUX21X1 U158 (rec_dataH_rec[5], rec_dataH_temp[4], test_se, n146);
  MUX21X1 U159 (n151, rec_dataH_rec[4], test_se, n147);
  MUX21X1 U160 (rec_dataH_temp[6], rec_dataH[5], test_se, n148);
  MUX21X1 U161 (rec_dataH_rec[6], rec_dataH_temp[5], test_se, n149);
  MUX21X1 U162 (n158, rec_dataH_rec[5], test_se, n150);
  MUX21X1 U163 (rec_dataH_temp[7], rec_dataH[6], test_se, n152);
  MUX21X1 U164 (rec_dataH_rec[7], rec_dataH_temp[6], test_se, n153);
  MUX21X1 U165 (n165, rec_dataH_rec[6], test_se, n154);
  MUX21X1 U166 (iRECEIVER_rec_readyInH, iRECEIVER_rec_datSyncH, test_se, n155);
wire iXMIT_xmit_doneInH (U213, U49);
wire iXMIT_next_state_0_ (U204, U110);
wire iXMIT_next_state_1_ (U207, U104);
wire iXMIT_next_state_2_ (U74, U105);
wire iXMIT_state_0_ (U97, U75, U71, U4, iXMIT_state_reg_0_, U104);
wire iXMIT_state_2_ (U83, U77, U71, U4, U3, iXMIT_state_reg_2_, U122);
wire iXMIT_bitCountH_0_ (U219, U208, U85, U65, iXMIT_bitCountH_reg_0_, U98);
wire iXMIT_bitCountH_1_ (U219, U208, U85, U63, iXMIT_bitCountH_reg_1_, U86);
wire iXMIT_bitCountH_2_ (U85, U61, iXMIT_bitCountH_reg_2_, U84);
wire iXMIT_bitCountH_3_ (U222, U59, iXMIT_bitCountH_reg_3_, U110);
wire iXMIT_N29 (U87, U134);
wire iXMIT_N28 (U294, U88, U115);
wire iXMIT_N27 (U294, U89, U130);
wire iXMIT_N26 (U294, U90, U133);
wire iXMIT_bitCell_cntrH_0_ (U215, U211, U94, iXMIT_bitCell_cntrH_reg_0_, U130);
wire iXMIT_bitCell_cntrH_1_ (U215, U211, U102, iXMIT_bitCell_cntrH_reg_1_, U115);
wire iXMIT_bitCell_cntrH_2_ (U102, iXMIT_bitCell_cntrH_reg_2_, U134);
wire iXMIT_bitCell_cntrH_3_ (U218, U102, iXMIT_bitCell_cntrH_reg_3_, U103);
wire iXMIT_xmit_ShiftRegH_1_ (U33, iXMIT_xmit_ShiftRegH_reg_1_, U53);
wire iXMIT_xmit_ShiftRegH_2_ (U36, iXMIT_xmit_ShiftRegH_reg_2_, U54);
wire iXMIT_xmit_ShiftRegH_3_ (U39, iXMIT_xmit_ShiftRegH_reg_3_, U70);
wire iXMIT_xmit_ShiftRegH_4_ (U42, iXMIT_xmit_ShiftRegH_reg_4_, U76);
wire iXMIT_xmit_ShiftRegH_5_ (U295, U45, iXMIT_xmit_ShiftRegH_reg_5_, U78);
wire iXMIT_xmit_ShiftRegH_6_ (U295, U48, iXMIT_xmit_ShiftRegH_reg_6_, U81);
wire iXMIT_xmit_ShiftRegH_7_ (U295, U56, U51, iXMIT_xmit_ShiftRegH_reg_7_, U49);
wire iRECEIVER_rec_readyInH (U106, U166);
wire iRECEIVER_next_state_0_ (U116, U43);
wire iRECEIVER_next_state_1_ (U109, U46);
wire iRECEIVER_next_state_2_ (U297, U108, U1);
wire iRECEIVER_state_0_ (U297, U135, U113, U111, iRECEIVER_state_reg_0_, U46);
wire iRECEIVER_state_1_ (U297, U117, U114, U15, iRECEIVER_state_reg_1_, U1);
wire iRECEIVER_state_2_ (U297, U129, iRECEIVER_state_reg_2_, U133);
wire iRECEIVER_recd_bitCntrH_0_ (U227, U210, U11, iRECEIVER_recd_bitCntrH_reg_0_, U139);
wire iRECEIVER_recd_bitCntrH_1_ (U227, U210, U120, U9, iRECEIVER_recd_bitCntrH_reg_1_, U136);
wire iRECEIVER_recd_bitCntrH_2_ (U120, U7, iRECEIVER_recd_bitCntrH_reg_2_, U141);
wire iRECEIVER_recd_bitCntrH_3_ (U230, U118, U13, iRECEIVER_recd_bitCntrH_reg_3_, U43);
wire iRECEIVER_N23 (U298, U124, U2);
wire iRECEIVER_N22 (U299, U125, U34);
wire iRECEIVER_N21 (U299, U126, U37);
wire iRECEIVER_N20 (U299, U127, U40);
wire iRECEIVER_bitCell_cntrH_0_ (U300, U223, U212, iRECEIVER_bitCell_cntrH_reg_0_, U37);
wire iRECEIVER_bitCell_cntrH_1_ (U300, U223, U212, U138, iRECEIVER_bitCell_cntrH_reg_1_, U34);
wire iRECEIVER_bitCell_cntrH_2_ (U138, U132, iRECEIVER_bitCell_cntrH_reg_2_, U2);
wire iRECEIVER_bitCell_cntrH_3_ (U226, U138, iRECEIVER_bitCell_cntrH_reg_3_, U144);
wire iRECEIVER_rec_datSyncH (iRECEIVER_rec_datSyncH_reg, U119, U166);
wire iRECEIVER_rec_datH (U117, U107, U31, iRECEIVER_rec_datH_reg, U121);
wire n100 (U6, U136);
wire n103 (U8, U139);
wire n106 (U10, U140);
wire n109 (U12, U141);
wire n116 (U16, U144);
wire n123 (U18, U147);
wire n130 (U20, U150);
wire n137 (U22, U153);
wire n144 (U24, U156);
wire n151 (U26, U159);
wire n158 (U28, U162);
wire n165 (U30, U165);
wire n190 (U32, U122);
wire n193 (U35, U52);
wire n196 (U38, U53);
wire n199 (U41, U54);
wire n202 (U44, U70);
wire n205 (U47, U76);
wire n208 (U50, U78);
wire n211 (U205, U81);
wire n214 (U58, U84);
wire n217 (U60, U86);
wire n220 (U62, U98);
wire n223 (U64, U103);
wire n238 (U116, U112, U111, U107, U106, U15, U14, iRECEIVER_state_reg_2_);
wire n239 (U293, U95, U91, U83, U77, U5, iXMIT_state_reg_0_);
wire n241 (U135, U123, U117, U112, U107, iRECEIVER_state_reg_1_);
wire n242 (U293, U100, U79, U72, U5, iXMIT_state_reg_2_);
wire n243 (U118, U11, iRECEIVER_recd_bitCntrH_reg_0_);
wire n244 (U132, iRECEIVER_bitCell_cntrH_reg_1_);
wire n245 (U129, U123, U106, U14, iRECEIVER_state_reg_0_);
wire n246 (U293, U97, U95, U79, U72, iXMIT_state_reg_1_);
wire n247 (U221, U220, iXMIT_bitCountH_reg_2_);
wire n248 (U114, U112, U15, iRECEIVER_rec_datH_reg);
wire n249 (U225, U224, iRECEIVER_bitCell_cntrH_reg_2_);
wire n250 (U229, U228, iRECEIVER_recd_bitCntrH_reg_2_);
wire n251 (U293, U217, U216, iXMIT_bitCell_cntrH_reg_2_);
wire n252 (U65, iXMIT_bitCountH_reg_0_);
wire n253 (U85, iXMIT_bitCountH_reg_3_);
wire n254 (U101, U90, iXMIT_bitCell_cntrH_reg_0_);
wire n255 (U138, U132, U127, iRECEIVER_bitCell_cntrH_reg_0_);
wire n256 (U132, iRECEIVER_bitCell_cntrH_reg_3_);
wire n257 (U32, U5, iXMIT_xmit_ShiftRegH_reg_0_);
wire n258 (U50, iXMIT_xmit_ShiftRegH_reg_6_);
wire n259 (U47, iXMIT_xmit_ShiftRegH_reg_5_);
wire n260 (U44, iXMIT_xmit_ShiftRegH_reg_4_);
wire n261 (U41, iXMIT_xmit_ShiftRegH_reg_3_);
wire n262 (U38, iXMIT_xmit_ShiftRegH_reg_2_);
wire n263 (U35, iXMIT_xmit_ShiftRegH_reg_1_);
wire test_pointTM (test_pointTM, U289);
wire n281 (iXMIT_xmit_ShiftRegH_reg_0_, U52);
wire xmit_doneH_temp (U303, iXMIT_xmit_doneH_reg, U142);
wire rec_dataH_rec_0_temp (U17, iRECEIVER_par_dataH_reg_0_, U143, U147);
wire iXMIT_state_1_temp (U305, U80, iXMIT_state_reg_1_, U105);
wire n94 (U129, U128);
wire n93 (U135, U128);
wire n92 (U128, U127, U126, U125, U124);
wire n91 (U201, U138, U137);
wire n9 (U201, U138, U137, U135, U129, U128, U127, U126, U125, U124, U14, U13, U11, U9, U7);
wire n89 (U120, U118);
wire n88 (U131, U129, U117);
wire n87 (U117, U116);
wire n86 (U118, U116);
wire n85 (U132, U131, U114);
wire n84 (U114, U113);
wire n83 (U201, U116, U109);
wire n82 (U112, U109);
wire n81 (U113, U109);
wire n80 (U201, U123, U118, U108);
wire n8 (U202, U201, U132, U131, U129, U123, U120, U118, U117, U116, U114, U113, U112, U111, U109, U108, U31, U29, U27, U25, U23, U21, U19, U17, U13, U11, U9, U7);
wire n79 (U137, U135, U108);
wire n77 (U107, U106);
wire n75 (U102, U101, U94);
wire n74 (U96, U92);
wire n73 (U92, U91);
wire n72 (U99, U91);
wire n71 (U91, U90, U89, U88, U87);
wire n7 (U137, U135, U108, U107, U106, U102, U101, U99, U96, U94, U92, U91, U90, U89, U88, U87, U7, U6);
wire n69 (U209, U85);
wire n68 (U204, U82);
wire n67 (U204, U83);
wire n66 (U97, U92, U82, U80);
wire n65 (U93, U92, U80);
wire n64 (U214, U79);
wire n63 (U207, U80);
wire n62 (U100, U99, U82, U75);
wire n61 (U209, U94, U93, U75);
wire n60 (U75, U74);
wire n58 (U73, U72);
wire n57 (U101, U100, U96, U82, U71);
wire n56 (U213, U71);
wire n55 (U213, U72, U69);
wire n54 (U95, U92, U83, U75, U68);
wire n53 (U209, U83, U67);
wire n52 (U68, U67);
wire n51 (U69, U66);
wire n50 (U65, U64);
wire n49 (U63, U62);
wire n48 (U61, U60);
wire n47 (U67, U66, U65, U63, U61, U59);
wire n46 (U66, U65, U63, U61, U59);
wire n45 (U59, U58);
wire n44 (U207, U77, U57, U56, U55);
wire n43 (U206, U205);
wire n42 (U205, U56);
wire n41 (U51, U50);
wire n39 (U48, U47);
wire n37 (U45, U44, U290, U289, U291);
wire n35 (U42, U41);
wire n33 (U39, U38);
wire n31 (U36, U35);
wire n3 (U48, U47, U45, U44, U42, U41, U39, U38, U36, U35, U5, U4, U290, U289, U291);
wire n29 (U57, U56, U51, U48, U45, U42, U39, U36, U33);
wire n28 (U214, U77, U57, U51, U48, U45, U42, U39, U36, U33, iXMIT_xmit_ShiftRegH_reg_0_, U52);
wire n275 (U230, U229);
wire n274 (U229, U228, U210);
wire n273 (U226, U225);
wire n272 (U225, U224, U212);
wire n271 (U222, U221);
wire n270 (U221, U220, U208);
wire n27 (U230, U229, U228, U226, U225, U224, U222, U221, U220, U212, U210, U208, U33, U32);
wire n269 (U218, U217);
wire n268 (U217, U216, U211);
wire n26 (U218, U217, U216, U211, U206, U55, U50, U47, U44, U41, U38, U35, U32, iXMIT_xmit_ShiftRegH_reg_4_, iXMIT_xmit_ShiftRegH_reg_3_, iXMIT_xmit_ShiftRegH_reg_2_, iXMIT_xmit_ShiftRegH_reg_1_);
wire n25 (U293, U229, U228, U217, U216, U138, U132, U127, U101, U90, U85, U65, U50, U47, U32, U31, U30, U5, iXMIT_bitCell_cntrH_reg_2_, iXMIT_bitCountH_reg_0_, iXMIT_bitCountH_reg_3_, iXMIT_xmit_ShiftRegH_reg_6_, iXMIT_xmit_ShiftRegH_reg_5_, iRECEIVER_bitCell_cntrH_reg_0_, iRECEIVER_bitCell_cntrH_reg_3_, iRECEIVER_recd_bitCntrH_reg_2_, iXMIT_bitCell_cntrH_reg_0_, iXMIT_xmit_ShiftRegH_reg_0_);
wire n24 (U293, U225, U224, U221, U220, U135, U132, U129, U123, U118, U117, U114, U112, U107, U106, U100, U97, U95, U79, U72, U29, U28, U15, U14, U11, U5, iXMIT_state_reg_2_, iXMIT_state_reg_1_, iXMIT_bitCountH_reg_2_, iRECEIVER_state_reg_1_, iRECEIVER_state_reg_0_, iRECEIVER_bitCell_cntrH_reg_1_, iRECEIVER_bitCell_cntrH_reg_2_, iRECEIVER_recd_bitCntrH_reg_0_, iRECEIVER_rec_datH_reg);
wire n23 (U293, U116, U112, U111, U107, U106, U95, U91, U83, U77, U27, U26, U15, U14, U5, iXMIT_state_reg_0_, iRECEIVER_state_reg_2_);
wire n22 (U64, U62, U25, U24, U98, U103);
wire n21 (U205, U60, U58, U23, U22, U81, U84, U86);
wire n20 (U50, U47, U44, U21, U20, U70, U76, U78);
wire n2 (U293, U230, U229, U228, U226, U225, U224, U222, U221, U220, U218, U217, U216, U214, U212, U211, U210, U208, U206, U205, U138, U135, U132, U129, U127, U123, U118, U117, U116, U114, U112, U111, U107, U106, U101, U100, U97, U95, U91, U90, U85, U83, U79, U77, U72, U65, U64, U62, U60, U58, U57, U56, U55, U51, U50, U48, U47, U45, U44, U42, U41, U39, U38, U36, U35, U33, U32, U31, U30, U29, U28, U27, U26, U25, U24, U23, U22, U21, U20, U15, U14, U11, U5, U4, U3, iXMIT_bitCell_cntrH_reg_2_, iXMIT_state_reg_0_, iXMIT_state_reg_2_, iXMIT_state_reg_1_, iXMIT_bitCountH_reg_0_, iXMIT_bitCountH_reg_2_, iXMIT_bitCountH_reg_3_, iXMIT_xmit_ShiftRegH_reg_6_, iXMIT_xmit_ShiftRegH_reg_5_, iXMIT_xmit_ShiftRegH_reg_4_, iXMIT_xmit_ShiftRegH_reg_3_, iXMIT_xmit_ShiftRegH_reg_2_, iXMIT_xmit_ShiftRegH_reg_1_, iRECEIVER_state_reg_1_, iRECEIVER_state_reg_0_, iRECEIVER_bitCell_cntrH_reg_0_, iRECEIVER_bitCell_cntrH_reg_1_, iRECEIVER_bitCell_cntrH_reg_2_, iRECEIVER_bitCell_cntrH_reg_3_, iRECEIVER_state_reg_2_, iRECEIVER_recd_bitCntrH_reg_0_, iRECEIVER_recd_bitCntrH_reg_2_, iXMIT_bitCell_cntrH_reg_0_, iXMIT_xmit_ShiftRegH_reg_0_, iRECEIVER_rec_datH_reg, U52, U70, U76, U78, U81, U84, U86, U98, U103);
wire n19 (U41, U38, U35, U32, U19, U18, U52, U53, U54, U122);
wire n18 (U202, U109, U31, U29, U27, U25, U23, U21, U19, U17, iXMIT_bitCell_cntrH_reg_2_, U115);
wire n17 (U17, U16, iXMIT_state_reg_0_, iXMIT_state_reg_2_, iXMIT_state_reg_1_, iXMIT_bitCountH_reg_0_, iXMIT_bitCountH_reg_1_, iXMIT_bitCountH_reg_2_, iXMIT_bitCountH_reg_3_, iXMIT_xmit_ShiftRegH_reg_7_, iXMIT_xmit_ShiftRegH_reg_6_, iXMIT_xmit_ShiftRegH_reg_5_, U76, U78, U81, U84, U86, U98, U103, U104, U105, U110);
wire n15 (U28, U26, U15, U14, iRECEIVER_bitCell_cntrH_reg_2_, iRECEIVER_bitCell_cntrH_reg_3_, iRECEIVER_state_reg_2_, iRECEIVER_rec_readyH_reg, iRECEIVER_par_dataH_reg_7_, rec_dataH_temp_reg_7_, rec_dataH_reg_7_, iRECEIVER_par_dataH_reg_6_, U1, U2, U34, U159, U162, U163, U164, U165, U166);
wire n12 (U18, U13, U12, iRECEIVER_par_dataH_reg_0_, rec_dataH_temp_reg_0_, rec_dataH_reg_0_, iRECEIVER_recd_bitCntrH_reg_3_, iRECEIVER_recd_bitCntrH_reg_0_, iRECEIVER_recd_bitCntrH_reg_1_, iRECEIVER_recd_bitCntrH_reg_2_, iXMIT_bitCell_cntrH_reg_3_, iXMIT_bitCell_cntrH_reg_0_, U133, U134, U136, U139, U140, U141, U142, U143, U144, U147);
wire n11 (U16, U11, U10, iXMIT_bitCell_cntrH_reg_1_, iXMIT_xmit_ShiftRegH_reg_0_, iRECEIVER_rec_datSyncH_reg, iRECEIVER_rec_datH_reg, U119, U121, U122, U130, U144);
wire n10 (U12, U10, U9, U8, U6, U136, U139, U140, U141);
wire iXMIT_xmit_CTRL (U296, U295);
wire iXMIT_state_1_ (U305, U80, U3, iXMIT_state_reg_1_, U105);
wire iXMIT_N_CTRL_2_ (U296, U294);
wire iXMIT_N_CTRL_1_ (U296, U293);
wire iXMIT_N46 (U222, U59);
wire iXMIT_N45 (U220, U61);
wire iXMIT_N44 (U219, U63);
wire iXMIT_N25 (U294, U218, U87);
wire iXMIT_N24 (U295, U216, U88);
wire iXMIT_N23 (U215, U89);
wire iXMIT_CRTL (U302, U296);
wire iRECEIVER_state_CTRL (U301, U297);
wire iRECEIVER_bitCell_CTRL (U301, U300);
wire iRECEIVER_N_CTRL_2_ (U301, U299);
wire iRECEIVER_N_CTRL_1_ (U301, U298);
wire iRECEIVER_N28 (U298, U230, U13);
wire iRECEIVER_N27 (U298, U228, U7);
wire iRECEIVER_N26 (U298, U227, U9);
wire iRECEIVER_N19 (U299, U226, U124);
wire iRECEIVER_N18 (U300, U224, U125);
wire iRECEIVER_N17 (U300, U223, U126);
wire iRECEIVER_CTRL (U302, U301);
wire iCTRL (U305, U303, U302);
wire test_pointDOUT (rec_dataH_temp_reg_7_, rec_dataH_temp_reg_6_, rec_dataH_temp_reg_5_, rec_dataH_temp_reg_4_, rec_dataH_temp_reg_3_, rec_dataH_temp_reg_2_, rec_dataH_temp_reg_1_, rec_dataH_temp_reg_0_, U291);
wire n371 (U290, U291);
wire n370 (U290, U289);
wire n115 (iRECEIVER_rec_datH_reg, U119);
wire n117 (iRECEIVER_rec_datSyncH_reg, U121);
wire n118 (iXMIT_xmit_ShiftRegH_reg_0_, U122);
wire n119 (iXMIT_bitCell_cntrH_reg_1_, U130);
wire n120 (iXMIT_bitCell_cntrH_reg_0_, U133);
wire n121 (iXMIT_bitCell_cntrH_reg_3_, U134);
wire n122 (iRECEIVER_recd_bitCntrH_reg_2_, U136);
wire n124 (iRECEIVER_recd_bitCntrH_reg_1_, U139);
wire n125 (iRECEIVER_recd_bitCntrH_reg_0_, U140);
wire n126 (iRECEIVER_recd_bitCntrH_reg_3_, U141);
wire n127 (rec_dataH_reg_0_, U142);
wire n128 (rec_dataH_temp_reg_0_, U143);
wire n129 (iRECEIVER_par_dataH_reg_0_, U144);
wire n131 (rec_dataH_reg_1_, U145);
wire n132 (rec_dataH_temp_reg_1_, U146);
wire n133 (iRECEIVER_par_dataH_reg_1_, U147);
wire n134 (rec_dataH_reg_2_, U148);
wire n135 (rec_dataH_temp_reg_2_, U149);
wire n136 (iRECEIVER_par_dataH_reg_2_, U150);
wire n138 (rec_dataH_reg_3_, U151);
wire n139 (rec_dataH_temp_reg_3_, U152);
wire n140 (iRECEIVER_par_dataH_reg_3_, U153);
wire n141 (rec_dataH_reg_4_, U154);
wire n142 (rec_dataH_temp_reg_4_, U155);
wire n143 (iRECEIVER_par_dataH_reg_4_, U156);
wire n145 (rec_dataH_reg_5_, U157);
wire n146 (rec_dataH_temp_reg_5_, U158);
wire n147 (iRECEIVER_par_dataH_reg_5_, U159);
wire n148 (rec_dataH_reg_6_, U160);
wire n149 (rec_dataH_temp_reg_6_, U161);
wire n150 (iRECEIVER_par_dataH_reg_6_, U162);
wire n152 (rec_dataH_reg_7_, U163);
wire n153 (rec_dataH_temp_reg_7_, U164);
wire n154 (iRECEIVER_par_dataH_reg_7_, U165);
wire n155 (iRECEIVER_rec_readyH_reg, U166);
wire n156 (iRECEIVER_state_reg_2_, U1);
wire n157 (iRECEIVER_bitCell_cntrH_reg_3_, U2);
wire n159 (iRECEIVER_bitCell_cntrH_reg_2_, U34);
wire n160 (iRECEIVER_bitCell_cntrH_reg_1_, U37);
wire n161 (iRECEIVER_bitCell_cntrH_reg_0_, U40);
wire n162 (iRECEIVER_state_reg_0_, U43);
wire n163 (iRECEIVER_state_reg_1_, U46);
wire n164 (iXMIT_xmit_doneH_reg, U49);
wire n166 (iXMIT_xmit_ShiftRegH_reg_1_, U52);
wire n167 (iXMIT_xmit_ShiftRegH_reg_2_, U53);
wire n168 (iXMIT_xmit_ShiftRegH_reg_3_, U54);
wire n169 (iXMIT_xmit_ShiftRegH_reg_4_, U70);
wire n170 (iXMIT_xmit_ShiftRegH_reg_5_, U76);
wire n171 (iXMIT_xmit_ShiftRegH_reg_6_, U78);
wire n172 (iXMIT_xmit_ShiftRegH_reg_7_, U81);
wire n173 (iXMIT_bitCountH_reg_3_, U84);
wire n174 (iXMIT_bitCountH_reg_2_, U86);
wire n175 (iXMIT_bitCountH_reg_1_, U98);
wire n176 (iXMIT_bitCountH_reg_0_, U103);
wire n177 (iXMIT_state_reg_1_, U104);
wire n178 (iXMIT_state_reg_2_, U105);
wire n179 (iXMIT_state_reg_0_, U110);
wire n180 (iXMIT_bitCell_cntrH_reg_2_, U115);
wire rec_dataH_rec_0 (U17, iRECEIVER_par_dataH_reg_0_, U143, U147);
endmodule